`timescale 1us/1ns

// Declares a module with no input and output prots (used for testbench/simulation)
module func_ex1 ();
	
	// This function returns the sum of 2x8bit numbers 
	// An internal variable with the same name as the function is 
	// created inside it and is used for returning the value 
	function [8:0] sum (input [7:0] a, input [7:0] b);
		begin 
			sum = a + b	// Since a and b are 8-bit, their sum can be up to 9 bits(510 max)
		end 
	endfunction 

	// Variables used for stimulus 
	reg [7:0] a, b;	// Declares two 8-bit registers and b to hold input values for testing the function

	initial begin 
		$monitor ($time, "a=%d, b=%d, sum=%d", a,b, sum(a,b));
		#1 a=1; b=9;
		#1 a=13; b=66;
		#1 a=255; b=1;
		#1 a=255; b=255;
	end 

endmodule
